package Defines;

typedef 12 CTRL_ADDR_WIDTH;
typedef 64 CTRL_DATA_WIDTH;
typedef 128 ST_DATA_WIDTH;
typedef 0 ST_USER_WIDTH;

typedef 3 NUM_LAYERS;
typedef 32 NUM_L0_STREAMS;
typedef 16 NUM_L1_STREAMS;
typedef 16 NUM_L2_STREAMS;
// typedef  1 NUM_L3_STREAMS;
// typedef TAdd#(TAdd#(TAdd#(NUM_L3_STREAMS, NUM_L2_STREAMS), NUM_L1_STREAMS), NUM_L0_STREAMS) NUM_STREAMS;
typedef TAdd#(TAdd#(NUM_L2_STREAMS, NUM_L1_STREAMS), NUM_L0_STREAMS) NUM_STREAMS;
// typedef TMax#(TMax#(TMax#(NUM_L3_STREAMS, NUM_L2_STREAMS), NUM_L1_STREAMS), NUM_L0_STREAMS) MAX_STREAMS_PER_LAYER;
typedef TMax#(TMax#(NUM_L2_STREAMS, NUM_L1_STREAMS), NUM_L0_STREAMS) MAX_STREAMS_PER_LAYER;
typedef 2048 L0_BRAM_SIZE_TOTAL;
typedef 2048 L1_BRAM_SIZE_TOTAL;
typedef 1024 L2_BRAM_SIZE_TOTAL;
// typedef   16 L3_BRAM_SIZE_TOTAL;
// typedef TMax#(TMax#(TMax#(L3_BRAM_SIZE_TOTAL, L2_BRAM_SIZE_TOTAL), L1_BRAM_SIZE_TOTAL), L0_BRAM_SIZE_TOTAL) MAX_BRAM_SIZE_TOTAL;
typedef TMax#(TMax#(L2_BRAM_SIZE_TOTAL, L1_BRAM_SIZE_TOTAL), L0_BRAM_SIZE_TOTAL) MAX_BRAM_SIZE_TOTAL;
typedef TDiv#(L0_BRAM_SIZE_TOTAL, NUM_L0_STREAMS) L0_BRAM_SIZE_PER_ENGINE;
typedef TDiv#(L1_BRAM_SIZE_TOTAL, NUM_L1_STREAMS) L1_BRAM_SIZE_PER_ENGINE;
typedef TDiv#(L2_BRAM_SIZE_TOTAL, NUM_L2_STREAMS) L2_BRAM_SIZE_PER_ENGINE;
// typedef TDiv#(L3_BRAM_SIZE_TOTAL, NUM_L3_STREAMS) L3_BRAM_SIZE_PER_ENGINE;
// typedef TMax#(TMax#(TMax#(L3_BRAM_SIZE_PER_ENGINE, L2_BRAM_SIZE_PER_ENGINE), L1_BRAM_SIZE_PER_ENGINE), L0_BRAM_SIZE_PER_ENGINE) MAX_BRAM_SIZE_PER_ENGINE;
typedef TMax#(TMax#(L2_BRAM_SIZE_PER_ENGINE, L1_BRAM_SIZE_PER_ENGINE), L0_BRAM_SIZE_PER_ENGINE) MAX_BRAM_SIZE_PER_ENGINE;
typedef TLog#(MAX_BRAM_SIZE_PER_ENGINE) BRAM_ADDR_WIDTH;
typedef TAdd#(TLog#(TMul#(NUM_STREAMS, MAX_BRAM_SIZE_PER_ENGINE)), 1) MEM_IFC_ADDR_WIDTH; // add one bit in case number of streams is not a power of 2
typedef TAdd#(MEM_IFC_ADDR_WIDTH, 4) MEM_AXI_ADDR_WIDTH;
typedef 128 BRAM_DATA_WIDTH;
typedef TDiv#(BRAM_DATA_WIDTH, 8) BRAM_BE_WIDTH;

// BRAM size in rows of 128 bit for each layer in total
// Integer numEngines[valueOf(NUM_LAYERS)] = {valueOf(NUM_L0_STREAMS), valueOf(NUM_L1_STREAMS), valueOf(NUM_L2_STREAMS), valueOf(NUM_L3_STREAMS)};
// Integer bramSizeTotal[valueOf(NUM_LAYERS)] = {valueOf(L0_BRAM_SIZE_TOTAL), valueOf(L1_BRAM_SIZE_TOTAL), valueOf(L2_BRAM_SIZE_TOTAL), valueOf(L3_BRAM_SIZE_TOTAL)};
// Integer bramSizePerEngine[valueOf(NUM_LAYERS)] = {valueOf(L0_BRAM_SIZE_PER_ENGINE), valueOf(L1_BRAM_SIZE_PER_ENGINE), valueOf(L2_BRAM_SIZE_PER_ENGINE), valueOf(L3_BRAM_SIZE_PER_ENGINE)};
Integer numEngines[valueOf(NUM_LAYERS)] = {valueOf(NUM_L0_STREAMS), valueOf(NUM_L1_STREAMS), valueOf(NUM_L2_STREAMS)};
Integer bramSizeTotal[valueOf(NUM_LAYERS)] = {valueOf(L0_BRAM_SIZE_TOTAL), valueOf(L1_BRAM_SIZE_TOTAL), valueOf(L2_BRAM_SIZE_TOTAL)};
Integer bramSizePerEngine[valueOf(NUM_LAYERS)] = {valueOf(L0_BRAM_SIZE_PER_ENGINE), valueOf(L1_BRAM_SIZE_PER_ENGINE), valueOf(L2_BRAM_SIZE_PER_ENGINE)};

endpackage : Defines
